`ifndef TYPEDEFS_SVH
`define TYPEDEFS_SVH

typedef bit [7:0] u8_t;
typedef u8_t byte_t;

`endif
