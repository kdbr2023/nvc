package nvc_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "base/typedefs.svh"
    `include "base/format.svh"
    `include "base/packet.svh"
//  `include "base/payload.svh"

    `include "policy/packet_printer.svh"
endpackage
